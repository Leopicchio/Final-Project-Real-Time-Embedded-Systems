// main_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module main_system (
		input  wire        audio_0_external_interface_ADCDAT,                //                  audio_0_external_interface.ADCDAT
		input  wire        audio_0_external_interface_ADCLRCK,               //                                            .ADCLRCK
		input  wire        audio_0_external_interface_BCLK,                  //                                            .BCLK
		output wire        audio_0_external_interface_DACDAT,                //                                            .DACDAT
		input  wire        audio_0_external_interface_DACLRCK,               //                                            .DACLRCK
		inout  wire        audio_and_video_config_0_external_interface_SDAT, // audio_and_video_config_0_external_interface.SDAT
		output wire        audio_and_video_config_0_external_interface_SCLK, //                                            .SCLK
		input  wire        clk_clk,                                          //                                         clk.clk
		output wire        clk_audio_codec_clk,                              //                             clk_audio_codec.clk
		output wire        clk_sdram_clk,                                    //                                   clk_sdram.clk
		input  wire [3:0]  pio_buttons_external_connection_export,           //             pio_buttons_external_connection.export
		output wire [9:0]  pio_leds_external_connection_export,              //                pio_leds_external_connection.export
		input  wire [9:0]  pio_switches_external_connection_export,          //            pio_switches_external_connection.export
		input  wire        reset_reset_n,                                    //                                       reset.reset_n
		output wire [12:0] sdram_controller_wire_addr,                       //                       sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,                         //                                            .ba
		output wire        sdram_controller_wire_cas_n,                      //                                            .cas_n
		output wire        sdram_controller_wire_cke,                        //                                            .cke
		output wire        sdram_controller_wire_cs_n,                       //                                            .cs_n
		inout  wire [15:0] sdram_controller_wire_dq,                         //                                            .dq
		output wire [1:0]  sdram_controller_wire_dqm,                        //                                            .dqm
		output wire        sdram_controller_wire_ras_n,                      //                                            .ras_n
		output wire        sdram_controller_wire_we_n,                       //                                            .we_n
		input  wire        uart_0_external_connection_rxd,                   //                  uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd                    //                                            .txd
	);

	wire         pll_outclk0_clk;                                                               // pll:outclk_0 -> [audio_0:clk, audio_and_video_config_0:clk, irq_mapper:clk, irq_mapper_001:clk, jtag_uart_0:clk, jtag_uart_1:clk, mailbox_simple_0:clk, mm_interconnect_0:pll_outclk0_clk, mutex_SDRAM:clk, nios2_FFT:clk, nios2_sound_acquisition:clk, onchip_memory:clk, onchip_memory_nios2_FFT:clk, pio_LEDS:clk, pio_buttons:clk, pio_switches:clk, rst_controller_001:clk, rst_controller_002:clk, sysid_qsys_0:clock, uart_0:clk]
	wire         pll_outclk1_clk;                                                               // pll:outclk_1 -> [SDRAM_controller:clk, mm_interconnect_0:pll_outclk1_clk, rst_controller:clk]
	wire  [31:0] nios2_sound_acquisition_data_master_readdata;                                  // mm_interconnect_0:nios2_sound_acquisition_data_master_readdata -> nios2_sound_acquisition:d_readdata
	wire         nios2_sound_acquisition_data_master_waitrequest;                               // mm_interconnect_0:nios2_sound_acquisition_data_master_waitrequest -> nios2_sound_acquisition:d_waitrequest
	wire         nios2_sound_acquisition_data_master_debugaccess;                               // nios2_sound_acquisition:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_sound_acquisition_data_master_debugaccess
	wire  [27:0] nios2_sound_acquisition_data_master_address;                                   // nios2_sound_acquisition:d_address -> mm_interconnect_0:nios2_sound_acquisition_data_master_address
	wire   [3:0] nios2_sound_acquisition_data_master_byteenable;                                // nios2_sound_acquisition:d_byteenable -> mm_interconnect_0:nios2_sound_acquisition_data_master_byteenable
	wire         nios2_sound_acquisition_data_master_read;                                      // nios2_sound_acquisition:d_read -> mm_interconnect_0:nios2_sound_acquisition_data_master_read
	wire         nios2_sound_acquisition_data_master_readdatavalid;                             // mm_interconnect_0:nios2_sound_acquisition_data_master_readdatavalid -> nios2_sound_acquisition:d_readdatavalid
	wire         nios2_sound_acquisition_data_master_write;                                     // nios2_sound_acquisition:d_write -> mm_interconnect_0:nios2_sound_acquisition_data_master_write
	wire  [31:0] nios2_sound_acquisition_data_master_writedata;                                 // nios2_sound_acquisition:d_writedata -> mm_interconnect_0:nios2_sound_acquisition_data_master_writedata
	wire  [31:0] nios2_fft_data_master_readdata;                                                // mm_interconnect_0:nios2_FFT_data_master_readdata -> nios2_FFT:d_readdata
	wire         nios2_fft_data_master_waitrequest;                                             // mm_interconnect_0:nios2_FFT_data_master_waitrequest -> nios2_FFT:d_waitrequest
	wire         nios2_fft_data_master_debugaccess;                                             // nios2_FFT:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_FFT_data_master_debugaccess
	wire  [27:0] nios2_fft_data_master_address;                                                 // nios2_FFT:d_address -> mm_interconnect_0:nios2_FFT_data_master_address
	wire   [3:0] nios2_fft_data_master_byteenable;                                              // nios2_FFT:d_byteenable -> mm_interconnect_0:nios2_FFT_data_master_byteenable
	wire         nios2_fft_data_master_read;                                                    // nios2_FFT:d_read -> mm_interconnect_0:nios2_FFT_data_master_read
	wire         nios2_fft_data_master_readdatavalid;                                           // mm_interconnect_0:nios2_FFT_data_master_readdatavalid -> nios2_FFT:d_readdatavalid
	wire         nios2_fft_data_master_write;                                                   // nios2_FFT:d_write -> mm_interconnect_0:nios2_FFT_data_master_write
	wire  [31:0] nios2_fft_data_master_writedata;                                               // nios2_FFT:d_writedata -> mm_interconnect_0:nios2_FFT_data_master_writedata
	wire  [31:0] nios2_fft_instruction_master_readdata;                                         // mm_interconnect_0:nios2_FFT_instruction_master_readdata -> nios2_FFT:i_readdata
	wire         nios2_fft_instruction_master_waitrequest;                                      // mm_interconnect_0:nios2_FFT_instruction_master_waitrequest -> nios2_FFT:i_waitrequest
	wire  [18:0] nios2_fft_instruction_master_address;                                          // nios2_FFT:i_address -> mm_interconnect_0:nios2_FFT_instruction_master_address
	wire         nios2_fft_instruction_master_read;                                             // nios2_FFT:i_read -> mm_interconnect_0:nios2_FFT_instruction_master_read
	wire         nios2_fft_instruction_master_readdatavalid;                                    // mm_interconnect_0:nios2_FFT_instruction_master_readdatavalid -> nios2_FFT:i_readdatavalid
	wire  [31:0] nios2_sound_acquisition_instruction_master_readdata;                           // mm_interconnect_0:nios2_sound_acquisition_instruction_master_readdata -> nios2_sound_acquisition:i_readdata
	wire         nios2_sound_acquisition_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_sound_acquisition_instruction_master_waitrequest -> nios2_sound_acquisition:i_waitrequest
	wire  [27:0] nios2_sound_acquisition_instruction_master_address;                            // nios2_sound_acquisition:i_address -> mm_interconnect_0:nios2_sound_acquisition_instruction_master_address
	wire         nios2_sound_acquisition_instruction_master_read;                               // nios2_sound_acquisition:i_read -> mm_interconnect_0:nios2_sound_acquisition_instruction_master_read
	wire         nios2_sound_acquisition_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_sound_acquisition_instruction_master_readdatavalid -> nios2_sound_acquisition:i_readdatavalid
	wire         mm_interconnect_0_audio_0_avalon_audio_slave_chipselect;                       // mm_interconnect_0:audio_0_avalon_audio_slave_chipselect -> audio_0:chipselect
	wire  [31:0] mm_interconnect_0_audio_0_avalon_audio_slave_readdata;                         // audio_0:readdata -> mm_interconnect_0:audio_0_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_0_avalon_audio_slave_address;                          // mm_interconnect_0:audio_0_avalon_audio_slave_address -> audio_0:address
	wire         mm_interconnect_0_audio_0_avalon_audio_slave_read;                             // mm_interconnect_0:audio_0_avalon_audio_slave_read -> audio_0:read
	wire         mm_interconnect_0_audio_0_avalon_audio_slave_write;                            // mm_interconnect_0:audio_0_avalon_audio_slave_write -> audio_0:write
	wire  [31:0] mm_interconnect_0_audio_0_avalon_audio_slave_writedata;                        // mm_interconnect_0:audio_0_avalon_audio_slave_writedata -> audio_0:writedata
	wire  [31:0] mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata;    // audio_and_video_config_0:readdata -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest; // audio_and_video_config_0:waitrequest -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address;     // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_address -> audio_and_video_config_0:address
	wire         mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read;        // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_read -> audio_and_video_config_0:read
	wire   [3:0] mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable;  // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_byteenable -> audio_and_video_config_0:byteenable
	wire         mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write;       // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_write -> audio_and_video_config_0:write
	wire  [31:0] mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata;   // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_writedata -> audio_and_video_config_0:writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                      // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                   // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata;                   // mailbox_simple_0:avmm_snd_readdata -> mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_readdata
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest;                // mailbox_simple_0:avmm_snd_waitrequest -> mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_waitrequest
	wire   [1:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address;                    // mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_address -> mailbox_simple_0:avmm_snd_address
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read;                       // mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_read -> mailbox_simple_0:avmm_snd_read
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write;                      // mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_write -> mailbox_simple_0:avmm_snd_write
	wire  [31:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata;                  // mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_writedata -> mailbox_simple_0:avmm_snd_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                         // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                          // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_readdata;            // nios2_sound_acquisition:debug_mem_slave_readdata -> mm_interconnect_0:nios2_sound_acquisition_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_waitrequest;         // nios2_sound_acquisition:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_sound_acquisition_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_debugaccess;         // mm_interconnect_0:nios2_sound_acquisition_debug_mem_slave_debugaccess -> nios2_sound_acquisition:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_address;             // mm_interconnect_0:nios2_sound_acquisition_debug_mem_slave_address -> nios2_sound_acquisition:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_read;                // mm_interconnect_0:nios2_sound_acquisition_debug_mem_slave_read -> nios2_sound_acquisition:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_byteenable;          // mm_interconnect_0:nios2_sound_acquisition_debug_mem_slave_byteenable -> nios2_sound_acquisition:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_write;               // mm_interconnect_0:nios2_sound_acquisition_debug_mem_slave_write -> nios2_sound_acquisition:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_writedata;           // mm_interconnect_0:nios2_sound_acquisition_debug_mem_slave_writedata -> nios2_sound_acquisition:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                                 // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                                   // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory_s1_address;                                    // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                                 // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                                      // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                                  // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                                      // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;                              // mm_interconnect_0:SDRAM_controller_s1_chipselect -> SDRAM_controller:az_cs
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_readdata;                                // SDRAM_controller:za_data -> mm_interconnect_0:SDRAM_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;                             // SDRAM_controller:za_waitrequest -> mm_interconnect_0:SDRAM_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;                                 // mm_interconnect_0:SDRAM_controller_s1_address -> SDRAM_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                                    // mm_interconnect_0:SDRAM_controller_s1_read -> SDRAM_controller:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_controller_s1_byteenable;                              // mm_interconnect_0:SDRAM_controller_s1_byteenable -> SDRAM_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;                           // SDRAM_controller:za_valid -> mm_interconnect_0:SDRAM_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;                                   // mm_interconnect_0:SDRAM_controller_s1_write -> SDRAM_controller:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_writedata;                               // mm_interconnect_0:SDRAM_controller_s1_writedata -> SDRAM_controller:az_data
	wire         mm_interconnect_0_pio_buttons_s1_chipselect;                                   // mm_interconnect_0:pio_buttons_s1_chipselect -> pio_buttons:chipselect
	wire  [31:0] mm_interconnect_0_pio_buttons_s1_readdata;                                     // pio_buttons:readdata -> mm_interconnect_0:pio_buttons_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_buttons_s1_address;                                      // mm_interconnect_0:pio_buttons_s1_address -> pio_buttons:address
	wire         mm_interconnect_0_pio_buttons_s1_write;                                        // mm_interconnect_0:pio_buttons_s1_write -> pio_buttons:write_n
	wire  [31:0] mm_interconnect_0_pio_buttons_s1_writedata;                                    // mm_interconnect_0:pio_buttons_s1_writedata -> pio_buttons:writedata
	wire         mm_interconnect_0_pio_leds_s1_chipselect;                                      // mm_interconnect_0:pio_LEDS_s1_chipselect -> pio_LEDS:chipselect
	wire  [31:0] mm_interconnect_0_pio_leds_s1_readdata;                                        // pio_LEDS:readdata -> mm_interconnect_0:pio_LEDS_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_leds_s1_address;                                         // mm_interconnect_0:pio_LEDS_s1_address -> pio_LEDS:address
	wire         mm_interconnect_0_pio_leds_s1_write;                                           // mm_interconnect_0:pio_LEDS_s1_write -> pio_LEDS:write_n
	wire  [31:0] mm_interconnect_0_pio_leds_s1_writedata;                                       // mm_interconnect_0:pio_LEDS_s1_writedata -> pio_LEDS:writedata
	wire         mm_interconnect_0_mutex_sdram_s1_chipselect;                                   // mm_interconnect_0:mutex_SDRAM_s1_chipselect -> mutex_SDRAM:chipselect
	wire  [31:0] mm_interconnect_0_mutex_sdram_s1_readdata;                                     // mutex_SDRAM:data_to_cpu -> mm_interconnect_0:mutex_SDRAM_s1_readdata
	wire   [0:0] mm_interconnect_0_mutex_sdram_s1_address;                                      // mm_interconnect_0:mutex_SDRAM_s1_address -> mutex_SDRAM:address
	wire         mm_interconnect_0_mutex_sdram_s1_read;                                         // mm_interconnect_0:mutex_SDRAM_s1_read -> mutex_SDRAM:read
	wire         mm_interconnect_0_mutex_sdram_s1_write;                                        // mm_interconnect_0:mutex_SDRAM_s1_write -> mutex_SDRAM:write
	wire  [31:0] mm_interconnect_0_mutex_sdram_s1_writedata;                                    // mm_interconnect_0:mutex_SDRAM_s1_writedata -> mutex_SDRAM:data_from_cpu
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect;                    // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_chipselect -> jtag_uart_1:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata;                      // jtag_uart_1:av_readdata -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest;                   // jtag_uart_1:av_waitrequest -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address;                       // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_address -> jtag_uart_1:av_address
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read;                          // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_read -> jtag_uart_1:av_read_n
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write;                         // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_write -> jtag_uart_1:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata;                     // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_writedata -> jtag_uart_1:av_writedata
	wire  [31:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata;                 // mailbox_simple_0:avmm_rcv_readdata -> mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_readdata
	wire   [1:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address;                  // mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_address -> mailbox_simple_0:avmm_rcv_address
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read;                     // mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_read -> mailbox_simple_0:avmm_rcv_read
	wire         mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write;                    // mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_write -> mailbox_simple_0:avmm_rcv_write
	wire  [31:0] mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata;                // mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_writedata -> mailbox_simple_0:avmm_rcv_writedata
	wire  [31:0] mm_interconnect_0_nios2_fft_debug_mem_slave_readdata;                          // nios2_FFT:debug_mem_slave_readdata -> mm_interconnect_0:nios2_FFT_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_fft_debug_mem_slave_waitrequest;                       // nios2_FFT:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_FFT_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_fft_debug_mem_slave_debugaccess;                       // mm_interconnect_0:nios2_FFT_debug_mem_slave_debugaccess -> nios2_FFT:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_fft_debug_mem_slave_address;                           // mm_interconnect_0:nios2_FFT_debug_mem_slave_address -> nios2_FFT:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_fft_debug_mem_slave_read;                              // mm_interconnect_0:nios2_FFT_debug_mem_slave_read -> nios2_FFT:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_fft_debug_mem_slave_byteenable;                        // mm_interconnect_0:nios2_FFT_debug_mem_slave_byteenable -> nios2_FFT:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_fft_debug_mem_slave_write;                             // mm_interconnect_0:nios2_FFT_debug_mem_slave_write -> nios2_FFT:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_fft_debug_mem_slave_writedata;                         // mm_interconnect_0:nios2_FFT_debug_mem_slave_writedata -> nios2_FFT:debug_mem_slave_writedata
	wire         mm_interconnect_0_pio_switches_s1_chipselect;                                  // mm_interconnect_0:pio_switches_s1_chipselect -> pio_switches:chipselect
	wire  [31:0] mm_interconnect_0_pio_switches_s1_readdata;                                    // pio_switches:readdata -> mm_interconnect_0:pio_switches_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_switches_s1_address;                                     // mm_interconnect_0:pio_switches_s1_address -> pio_switches:address
	wire         mm_interconnect_0_pio_switches_s1_write;                                       // mm_interconnect_0:pio_switches_s1_write -> pio_switches:write_n
	wire  [31:0] mm_interconnect_0_pio_switches_s1_writedata;                                   // mm_interconnect_0:pio_switches_s1_writedata -> pio_switches:writedata
	wire         mm_interconnect_0_onchip_memory_nios2_fft_s1_chipselect;                       // mm_interconnect_0:onchip_memory_nios2_FFT_s1_chipselect -> onchip_memory_nios2_FFT:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_nios2_fft_s1_readdata;                         // onchip_memory_nios2_FFT:readdata -> mm_interconnect_0:onchip_memory_nios2_FFT_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory_nios2_fft_s1_address;                          // mm_interconnect_0:onchip_memory_nios2_FFT_s1_address -> onchip_memory_nios2_FFT:address
	wire   [3:0] mm_interconnect_0_onchip_memory_nios2_fft_s1_byteenable;                       // mm_interconnect_0:onchip_memory_nios2_FFT_s1_byteenable -> onchip_memory_nios2_FFT:byteenable
	wire         mm_interconnect_0_onchip_memory_nios2_fft_s1_write;                            // mm_interconnect_0:onchip_memory_nios2_FFT_s1_write -> onchip_memory_nios2_FFT:write
	wire  [31:0] mm_interconnect_0_onchip_memory_nios2_fft_s1_writedata;                        // mm_interconnect_0:onchip_memory_nios2_FFT_s1_writedata -> onchip_memory_nios2_FFT:writedata
	wire         mm_interconnect_0_onchip_memory_nios2_fft_s1_clken;                            // mm_interconnect_0:onchip_memory_nios2_FFT_s1_clken -> onchip_memory_nios2_FFT:clken
	wire         mm_interconnect_0_uart_0_s1_chipselect;                                        // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                                          // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                                           // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                              // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                                     // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                             // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                                         // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         irq_mapper_receiver0_irq;                                                      // mailbox_simple_0:irq_msg -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                      // uart_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                      // jtag_uart_1:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_fft_irq_irq;                                                             // irq_mapper:sender_irq -> nios2_FFT:irq
	wire         irq_mapper_001_receiver0_irq;                                                  // audio_0:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                                  // jtag_uart_0:av_irq -> irq_mapper_001:receiver1_irq
	wire         irq_mapper_001_receiver2_irq;                                                  // pio_buttons:irq -> irq_mapper_001:receiver2_irq
	wire  [31:0] nios2_sound_acquisition_irq_irq;                                               // irq_mapper_001:sender_irq -> nios2_sound_acquisition:irq
	wire         rst_controller_reset_out_reset;                                                // rst_controller:reset_out -> [SDRAM_controller:reset_n, mm_interconnect_0:SDRAM_controller_reset_reset_bridge_in_reset_reset]
	wire         nios2_sound_acquisition_debug_reset_request_reset;                             // nios2_sound_acquisition:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_003:reset_in1]
	wire         nios2_fft_debug_reset_request_reset;                                           // nios2_FFT:debug_reset_request -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in1, rst_controller_003:reset_in2]
	wire         rst_controller_001_reset_out_reset;                                            // rst_controller_001:reset_out -> [audio_0:reset, audio_and_video_config_0:reset, irq_mapper:reset, irq_mapper_001:reset, jtag_uart_0:rst_n, mailbox_simple_0:rst_n, mm_interconnect_0:nios2_sound_acquisition_reset_reset_bridge_in_reset_reset, mutex_SDRAM:reset_n, nios2_FFT:reset_n, nios2_sound_acquisition:reset_n, onchip_memory:reset, onchip_memory_nios2_FFT:reset, pio_LEDS:reset_n, pio_buttons:reset_n, pio_switches:reset_n, rst_translator:in_reset, sysid_qsys_0:reset_n, uart_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                                        // rst_controller_001:reset_req -> [nios2_FFT:reset_req, nios2_sound_acquisition:reset_req, onchip_memory:reset_req, onchip_memory_nios2_FFT:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                                            // rst_controller_002:reset_out -> [jtag_uart_1:rst_n, mm_interconnect_0:jtag_uart_1_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                                            // rst_controller_003:reset_out -> pll:rst

	main_system_SDRAM_controller sdram_controller (
		.clk            (pll_outclk1_clk),                                     //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                           //      .export
	);

	main_system_audio_0 audio_0 (
		.clk         (pll_outclk0_clk),                                         //                clk.clk
		.reset       (rst_controller_001_reset_out_reset),                      //              reset.reset
		.address     (mm_interconnect_0_audio_0_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_0_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_0_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_0_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_0_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_0_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_001_receiver0_irq),                            //          interrupt.irq
		.AUD_ADCDAT  (audio_0_external_interface_ADCDAT),                       // external_interface.export
		.AUD_ADCLRCK (audio_0_external_interface_ADCLRCK),                      //                   .export
		.AUD_BCLK    (audio_0_external_interface_BCLK),                         //                   .export
		.AUD_DACDAT  (audio_0_external_interface_DACDAT),                       //                   .export
		.AUD_DACLRCK (audio_0_external_interface_DACLRCK)                       //                   .export
	);

	main_system_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (pll_outclk0_clk),                                                               //                    clk.clk
		.reset       (rst_controller_001_reset_out_reset),                                            //                  reset.reset
		.address     (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_0_external_interface_SDAT),                              //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_0_external_interface_SCLK)                               //                       .export
	);

	main_system_jtag_uart_0 jtag_uart_0 (
		.clk            (pll_outclk0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                 //               irq.irq
	);

	main_system_jtag_uart_0 jtag_uart_1 (
		.clk            (pll_outclk0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                     //               irq.irq
	);

	altera_avalon_mailbox #(
		.DWIDTH (32),
		.AWIDTH (2)
	) mailbox_simple_0 (
		.clk                  (pll_outclk0_clk),                                                //                   clk.clk
		.rst_n                (~rst_controller_001_reset_out_reset),                            //                 rst_n.reset_n
		.avmm_snd_address     (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address),     //       avmm_msg_sender.address
		.avmm_snd_writedata   (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata),   //                      .writedata
		.avmm_snd_write       (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write),       //                      .write
		.avmm_snd_read        (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read),        //                      .read
		.avmm_snd_readdata    (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata),    //                      .readdata
		.avmm_snd_waitrequest (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest), //                      .waitrequest
		.irq_msg              (irq_mapper_receiver0_irq),                                       // interrupt_msg_pending.irq
		.avmm_rcv_address     (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address),   //     avmm_msg_receiver.address
		.avmm_rcv_read        (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read),      //                      .read
		.avmm_rcv_writedata   (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata), //                      .writedata
		.avmm_rcv_write       (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write),     //                      .write
		.avmm_rcv_readdata    (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata),  //                      .readdata
		.irq_space            ()                                                                //           (terminated)
	);

	main_system_mutex_SDRAM mutex_sdram (
		.reset_n       (~rst_controller_001_reset_out_reset),         // reset.reset_n
		.clk           (pll_outclk0_clk),                             //   clk.clk
		.chipselect    (mm_interconnect_0_mutex_sdram_s1_chipselect), //    s1.chipselect
		.data_from_cpu (mm_interconnect_0_mutex_sdram_s1_writedata),  //      .writedata
		.read          (mm_interconnect_0_mutex_sdram_s1_read),       //      .read
		.write         (mm_interconnect_0_mutex_sdram_s1_write),      //      .write
		.data_to_cpu   (mm_interconnect_0_mutex_sdram_s1_readdata),   //      .readdata
		.address       (mm_interconnect_0_mutex_sdram_s1_address)     //      .address
	);

	main_system_nios2_FFT nios2_fft (
		.clk                                 (pll_outclk0_clk),                                         //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_fft_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_fft_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_fft_data_master_read),                              //                          .read
		.d_readdata                          (nios2_fft_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_fft_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_fft_data_master_write),                             //                          .write
		.d_writedata                         (nios2_fft_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_fft_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_fft_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_fft_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_fft_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_fft_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_fft_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_fft_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_fft_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_fft_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_fft_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_fft_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_fft_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_fft_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_fft_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_fft_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_fft_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_fft_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	main_system_nios2_sound_acquisition nios2_sound_acquisition (
		.clk                                 (pll_outclk0_clk),                                                       //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                                   //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                                //                          .reset_req
		.d_address                           (nios2_sound_acquisition_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_sound_acquisition_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_sound_acquisition_data_master_read),                              //                          .read
		.d_readdata                          (nios2_sound_acquisition_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_sound_acquisition_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_sound_acquisition_data_master_write),                             //                          .write
		.d_writedata                         (nios2_sound_acquisition_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_sound_acquisition_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_sound_acquisition_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_sound_acquisition_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_sound_acquisition_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_sound_acquisition_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_sound_acquisition_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_sound_acquisition_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_sound_acquisition_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_sound_acquisition_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                                       // custom_instruction_master.readra
	);

	main_system_onchip_memory onchip_memory (
		.clk        (pll_outclk0_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),        //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	main_system_onchip_memory_nios2_FFT onchip_memory_nios2_fft (
		.clk        (pll_outclk0_clk),                                         //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_nios2_fft_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_nios2_fft_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_nios2_fft_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_nios2_fft_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_nios2_fft_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_nios2_fft_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_nios2_fft_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),                      // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),                  //       .reset_req
		.freeze     (1'b0)                                                     // (terminated)
	);

	main_system_pio_LEDS pio_leds (
		.clk        (pll_outclk0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_pio_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_leds_s1_readdata),   //                    .readdata
		.out_port   (pio_leds_external_connection_export)       // external_connection.export
	);

	main_system_pio_buttons pio_buttons (
		.clk        (pll_outclk0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_buttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_buttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_buttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_buttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_buttons_s1_readdata),   //                    .readdata
		.in_port    (pio_buttons_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver2_irq)                 //                 irq.irq
	);

	main_system_pio_switches pio_switches (
		.clk        (pll_outclk0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_pio_switches_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_switches_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_switches_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_switches_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_switches_s1_readdata),   //                    .readdata
		.in_port    (pio_switches_external_connection_export),      // external_connection.export
		.irq        ()                                              //                 irq.irq
	);

	main_system_pll pll (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_003_reset_out_reset), //   reset.reset
		.outclk_0 (pll_outclk0_clk),                    // outclk0.clk
		.outclk_1 (pll_outclk1_clk),                    // outclk1.clk
		.outclk_2 (clk_sdram_clk),                      // outclk2.clk
		.outclk_3 (clk_audio_codec_clk),                // outclk3.clk
		.locked   ()                                    // (terminated)
	);

	main_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (pll_outclk0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	main_system_uart_0 uart_0 (
		.clk           (pll_outclk0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver1_irq)                   //                 irq.irq
	);

	main_system_mm_interconnect_0 mm_interconnect_0 (
		.pll_outclk0_clk                                             (pll_outclk0_clk),                                                               //                                         pll_outclk0.clk
		.pll_outclk1_clk                                             (pll_outclk1_clk),                                                               //                                         pll_outclk1.clk
		.jtag_uart_1_reset_reset_bridge_in_reset_reset               (rst_controller_002_reset_out_reset),                                            //             jtag_uart_1_reset_reset_bridge_in_reset.reset
		.nios2_sound_acquisition_reset_reset_bridge_in_reset_reset   (rst_controller_001_reset_out_reset),                                            // nios2_sound_acquisition_reset_reset_bridge_in_reset.reset
		.SDRAM_controller_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                                                //        SDRAM_controller_reset_reset_bridge_in_reset.reset
		.nios2_FFT_data_master_address                               (nios2_fft_data_master_address),                                                 //                               nios2_FFT_data_master.address
		.nios2_FFT_data_master_waitrequest                           (nios2_fft_data_master_waitrequest),                                             //                                                    .waitrequest
		.nios2_FFT_data_master_byteenable                            (nios2_fft_data_master_byteenable),                                              //                                                    .byteenable
		.nios2_FFT_data_master_read                                  (nios2_fft_data_master_read),                                                    //                                                    .read
		.nios2_FFT_data_master_readdata                              (nios2_fft_data_master_readdata),                                                //                                                    .readdata
		.nios2_FFT_data_master_readdatavalid                         (nios2_fft_data_master_readdatavalid),                                           //                                                    .readdatavalid
		.nios2_FFT_data_master_write                                 (nios2_fft_data_master_write),                                                   //                                                    .write
		.nios2_FFT_data_master_writedata                             (nios2_fft_data_master_writedata),                                               //                                                    .writedata
		.nios2_FFT_data_master_debugaccess                           (nios2_fft_data_master_debugaccess),                                             //                                                    .debugaccess
		.nios2_FFT_instruction_master_address                        (nios2_fft_instruction_master_address),                                          //                        nios2_FFT_instruction_master.address
		.nios2_FFT_instruction_master_waitrequest                    (nios2_fft_instruction_master_waitrequest),                                      //                                                    .waitrequest
		.nios2_FFT_instruction_master_read                           (nios2_fft_instruction_master_read),                                             //                                                    .read
		.nios2_FFT_instruction_master_readdata                       (nios2_fft_instruction_master_readdata),                                         //                                                    .readdata
		.nios2_FFT_instruction_master_readdatavalid                  (nios2_fft_instruction_master_readdatavalid),                                    //                                                    .readdatavalid
		.nios2_sound_acquisition_data_master_address                 (nios2_sound_acquisition_data_master_address),                                   //                 nios2_sound_acquisition_data_master.address
		.nios2_sound_acquisition_data_master_waitrequest             (nios2_sound_acquisition_data_master_waitrequest),                               //                                                    .waitrequest
		.nios2_sound_acquisition_data_master_byteenable              (nios2_sound_acquisition_data_master_byteenable),                                //                                                    .byteenable
		.nios2_sound_acquisition_data_master_read                    (nios2_sound_acquisition_data_master_read),                                      //                                                    .read
		.nios2_sound_acquisition_data_master_readdata                (nios2_sound_acquisition_data_master_readdata),                                  //                                                    .readdata
		.nios2_sound_acquisition_data_master_readdatavalid           (nios2_sound_acquisition_data_master_readdatavalid),                             //                                                    .readdatavalid
		.nios2_sound_acquisition_data_master_write                   (nios2_sound_acquisition_data_master_write),                                     //                                                    .write
		.nios2_sound_acquisition_data_master_writedata               (nios2_sound_acquisition_data_master_writedata),                                 //                                                    .writedata
		.nios2_sound_acquisition_data_master_debugaccess             (nios2_sound_acquisition_data_master_debugaccess),                               //                                                    .debugaccess
		.nios2_sound_acquisition_instruction_master_address          (nios2_sound_acquisition_instruction_master_address),                            //          nios2_sound_acquisition_instruction_master.address
		.nios2_sound_acquisition_instruction_master_waitrequest      (nios2_sound_acquisition_instruction_master_waitrequest),                        //                                                    .waitrequest
		.nios2_sound_acquisition_instruction_master_read             (nios2_sound_acquisition_instruction_master_read),                               //                                                    .read
		.nios2_sound_acquisition_instruction_master_readdata         (nios2_sound_acquisition_instruction_master_readdata),                           //                                                    .readdata
		.nios2_sound_acquisition_instruction_master_readdatavalid    (nios2_sound_acquisition_instruction_master_readdatavalid),                      //                                                    .readdatavalid
		.audio_0_avalon_audio_slave_address                          (mm_interconnect_0_audio_0_avalon_audio_slave_address),                          //                          audio_0_avalon_audio_slave.address
		.audio_0_avalon_audio_slave_write                            (mm_interconnect_0_audio_0_avalon_audio_slave_write),                            //                                                    .write
		.audio_0_avalon_audio_slave_read                             (mm_interconnect_0_audio_0_avalon_audio_slave_read),                             //                                                    .read
		.audio_0_avalon_audio_slave_readdata                         (mm_interconnect_0_audio_0_avalon_audio_slave_readdata),                         //                                                    .readdata
		.audio_0_avalon_audio_slave_writedata                        (mm_interconnect_0_audio_0_avalon_audio_slave_writedata),                        //                                                    .writedata
		.audio_0_avalon_audio_slave_chipselect                       (mm_interconnect_0_audio_0_avalon_audio_slave_chipselect),                       //                                                    .chipselect
		.audio_and_video_config_0_avalon_av_config_slave_address     (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address),     //     audio_and_video_config_0_avalon_av_config_slave.address
		.audio_and_video_config_0_avalon_av_config_slave_write       (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write),       //                                                    .write
		.audio_and_video_config_0_avalon_av_config_slave_read        (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read),        //                                                    .read
		.audio_and_video_config_0_avalon_av_config_slave_readdata    (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata),    //                                                    .readdata
		.audio_and_video_config_0_avalon_av_config_slave_writedata   (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata),   //                                                    .writedata
		.audio_and_video_config_0_avalon_av_config_slave_byteenable  (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable),  //                                                    .byteenable
		.audio_and_video_config_0_avalon_av_config_slave_waitrequest (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest), //                                                    .waitrequest
		.jtag_uart_0_avalon_jtag_slave_address                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                       //                       jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                         //                                                    .write
		.jtag_uart_0_avalon_jtag_slave_read                          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                          //                                                    .read
		.jtag_uart_0_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                      //                                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                     //                                                    .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                   //                                                    .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                    //                                                    .chipselect
		.jtag_uart_1_avalon_jtag_slave_address                       (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),                       //                       jtag_uart_1_avalon_jtag_slave.address
		.jtag_uart_1_avalon_jtag_slave_write                         (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),                         //                                                    .write
		.jtag_uart_1_avalon_jtag_slave_read                          (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),                          //                                                    .read
		.jtag_uart_1_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),                      //                                                    .readdata
		.jtag_uart_1_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),                     //                                                    .writedata
		.jtag_uart_1_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest),                   //                                                    .waitrequest
		.jtag_uart_1_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),                    //                                                    .chipselect
		.mailbox_simple_0_avmm_msg_receiver_address                  (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address),                  //                  mailbox_simple_0_avmm_msg_receiver.address
		.mailbox_simple_0_avmm_msg_receiver_write                    (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write),                    //                                                    .write
		.mailbox_simple_0_avmm_msg_receiver_read                     (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read),                     //                                                    .read
		.mailbox_simple_0_avmm_msg_receiver_readdata                 (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata),                 //                                                    .readdata
		.mailbox_simple_0_avmm_msg_receiver_writedata                (mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata),                //                                                    .writedata
		.mailbox_simple_0_avmm_msg_sender_address                    (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address),                    //                    mailbox_simple_0_avmm_msg_sender.address
		.mailbox_simple_0_avmm_msg_sender_write                      (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write),                      //                                                    .write
		.mailbox_simple_0_avmm_msg_sender_read                       (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read),                       //                                                    .read
		.mailbox_simple_0_avmm_msg_sender_readdata                   (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata),                   //                                                    .readdata
		.mailbox_simple_0_avmm_msg_sender_writedata                  (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata),                  //                                                    .writedata
		.mailbox_simple_0_avmm_msg_sender_waitrequest                (mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest),                //                                                    .waitrequest
		.mutex_SDRAM_s1_address                                      (mm_interconnect_0_mutex_sdram_s1_address),                                      //                                      mutex_SDRAM_s1.address
		.mutex_SDRAM_s1_write                                        (mm_interconnect_0_mutex_sdram_s1_write),                                        //                                                    .write
		.mutex_SDRAM_s1_read                                         (mm_interconnect_0_mutex_sdram_s1_read),                                         //                                                    .read
		.mutex_SDRAM_s1_readdata                                     (mm_interconnect_0_mutex_sdram_s1_readdata),                                     //                                                    .readdata
		.mutex_SDRAM_s1_writedata                                    (mm_interconnect_0_mutex_sdram_s1_writedata),                                    //                                                    .writedata
		.mutex_SDRAM_s1_chipselect                                   (mm_interconnect_0_mutex_sdram_s1_chipselect),                                   //                                                    .chipselect
		.nios2_FFT_debug_mem_slave_address                           (mm_interconnect_0_nios2_fft_debug_mem_slave_address),                           //                           nios2_FFT_debug_mem_slave.address
		.nios2_FFT_debug_mem_slave_write                             (mm_interconnect_0_nios2_fft_debug_mem_slave_write),                             //                                                    .write
		.nios2_FFT_debug_mem_slave_read                              (mm_interconnect_0_nios2_fft_debug_mem_slave_read),                              //                                                    .read
		.nios2_FFT_debug_mem_slave_readdata                          (mm_interconnect_0_nios2_fft_debug_mem_slave_readdata),                          //                                                    .readdata
		.nios2_FFT_debug_mem_slave_writedata                         (mm_interconnect_0_nios2_fft_debug_mem_slave_writedata),                         //                                                    .writedata
		.nios2_FFT_debug_mem_slave_byteenable                        (mm_interconnect_0_nios2_fft_debug_mem_slave_byteenable),                        //                                                    .byteenable
		.nios2_FFT_debug_mem_slave_waitrequest                       (mm_interconnect_0_nios2_fft_debug_mem_slave_waitrequest),                       //                                                    .waitrequest
		.nios2_FFT_debug_mem_slave_debugaccess                       (mm_interconnect_0_nios2_fft_debug_mem_slave_debugaccess),                       //                                                    .debugaccess
		.nios2_sound_acquisition_debug_mem_slave_address             (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_address),             //             nios2_sound_acquisition_debug_mem_slave.address
		.nios2_sound_acquisition_debug_mem_slave_write               (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_write),               //                                                    .write
		.nios2_sound_acquisition_debug_mem_slave_read                (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_read),                //                                                    .read
		.nios2_sound_acquisition_debug_mem_slave_readdata            (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_readdata),            //                                                    .readdata
		.nios2_sound_acquisition_debug_mem_slave_writedata           (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_writedata),           //                                                    .writedata
		.nios2_sound_acquisition_debug_mem_slave_byteenable          (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_byteenable),          //                                                    .byteenable
		.nios2_sound_acquisition_debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_waitrequest),         //                                                    .waitrequest
		.nios2_sound_acquisition_debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_sound_acquisition_debug_mem_slave_debugaccess),         //                                                    .debugaccess
		.onchip_memory_s1_address                                    (mm_interconnect_0_onchip_memory_s1_address),                                    //                                    onchip_memory_s1.address
		.onchip_memory_s1_write                                      (mm_interconnect_0_onchip_memory_s1_write),                                      //                                                    .write
		.onchip_memory_s1_readdata                                   (mm_interconnect_0_onchip_memory_s1_readdata),                                   //                                                    .readdata
		.onchip_memory_s1_writedata                                  (mm_interconnect_0_onchip_memory_s1_writedata),                                  //                                                    .writedata
		.onchip_memory_s1_byteenable                                 (mm_interconnect_0_onchip_memory_s1_byteenable),                                 //                                                    .byteenable
		.onchip_memory_s1_chipselect                                 (mm_interconnect_0_onchip_memory_s1_chipselect),                                 //                                                    .chipselect
		.onchip_memory_s1_clken                                      (mm_interconnect_0_onchip_memory_s1_clken),                                      //                                                    .clken
		.onchip_memory_nios2_FFT_s1_address                          (mm_interconnect_0_onchip_memory_nios2_fft_s1_address),                          //                          onchip_memory_nios2_FFT_s1.address
		.onchip_memory_nios2_FFT_s1_write                            (mm_interconnect_0_onchip_memory_nios2_fft_s1_write),                            //                                                    .write
		.onchip_memory_nios2_FFT_s1_readdata                         (mm_interconnect_0_onchip_memory_nios2_fft_s1_readdata),                         //                                                    .readdata
		.onchip_memory_nios2_FFT_s1_writedata                        (mm_interconnect_0_onchip_memory_nios2_fft_s1_writedata),                        //                                                    .writedata
		.onchip_memory_nios2_FFT_s1_byteenable                       (mm_interconnect_0_onchip_memory_nios2_fft_s1_byteenable),                       //                                                    .byteenable
		.onchip_memory_nios2_FFT_s1_chipselect                       (mm_interconnect_0_onchip_memory_nios2_fft_s1_chipselect),                       //                                                    .chipselect
		.onchip_memory_nios2_FFT_s1_clken                            (mm_interconnect_0_onchip_memory_nios2_fft_s1_clken),                            //                                                    .clken
		.pio_buttons_s1_address                                      (mm_interconnect_0_pio_buttons_s1_address),                                      //                                      pio_buttons_s1.address
		.pio_buttons_s1_write                                        (mm_interconnect_0_pio_buttons_s1_write),                                        //                                                    .write
		.pio_buttons_s1_readdata                                     (mm_interconnect_0_pio_buttons_s1_readdata),                                     //                                                    .readdata
		.pio_buttons_s1_writedata                                    (mm_interconnect_0_pio_buttons_s1_writedata),                                    //                                                    .writedata
		.pio_buttons_s1_chipselect                                   (mm_interconnect_0_pio_buttons_s1_chipselect),                                   //                                                    .chipselect
		.pio_LEDS_s1_address                                         (mm_interconnect_0_pio_leds_s1_address),                                         //                                         pio_LEDS_s1.address
		.pio_LEDS_s1_write                                           (mm_interconnect_0_pio_leds_s1_write),                                           //                                                    .write
		.pio_LEDS_s1_readdata                                        (mm_interconnect_0_pio_leds_s1_readdata),                                        //                                                    .readdata
		.pio_LEDS_s1_writedata                                       (mm_interconnect_0_pio_leds_s1_writedata),                                       //                                                    .writedata
		.pio_LEDS_s1_chipselect                                      (mm_interconnect_0_pio_leds_s1_chipselect),                                      //                                                    .chipselect
		.pio_switches_s1_address                                     (mm_interconnect_0_pio_switches_s1_address),                                     //                                     pio_switches_s1.address
		.pio_switches_s1_write                                       (mm_interconnect_0_pio_switches_s1_write),                                       //                                                    .write
		.pio_switches_s1_readdata                                    (mm_interconnect_0_pio_switches_s1_readdata),                                    //                                                    .readdata
		.pio_switches_s1_writedata                                   (mm_interconnect_0_pio_switches_s1_writedata),                                   //                                                    .writedata
		.pio_switches_s1_chipselect                                  (mm_interconnect_0_pio_switches_s1_chipselect),                                  //                                                    .chipselect
		.SDRAM_controller_s1_address                                 (mm_interconnect_0_sdram_controller_s1_address),                                 //                                 SDRAM_controller_s1.address
		.SDRAM_controller_s1_write                                   (mm_interconnect_0_sdram_controller_s1_write),                                   //                                                    .write
		.SDRAM_controller_s1_read                                    (mm_interconnect_0_sdram_controller_s1_read),                                    //                                                    .read
		.SDRAM_controller_s1_readdata                                (mm_interconnect_0_sdram_controller_s1_readdata),                                //                                                    .readdata
		.SDRAM_controller_s1_writedata                               (mm_interconnect_0_sdram_controller_s1_writedata),                               //                                                    .writedata
		.SDRAM_controller_s1_byteenable                              (mm_interconnect_0_sdram_controller_s1_byteenable),                              //                                                    .byteenable
		.SDRAM_controller_s1_readdatavalid                           (mm_interconnect_0_sdram_controller_s1_readdatavalid),                           //                                                    .readdatavalid
		.SDRAM_controller_s1_waitrequest                             (mm_interconnect_0_sdram_controller_s1_waitrequest),                             //                                                    .waitrequest
		.SDRAM_controller_s1_chipselect                              (mm_interconnect_0_sdram_controller_s1_chipselect),                              //                                                    .chipselect
		.sysid_qsys_0_control_slave_address                          (mm_interconnect_0_sysid_qsys_0_control_slave_address),                          //                          sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                         (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                         //                                                    .readdata
		.uart_0_s1_address                                           (mm_interconnect_0_uart_0_s1_address),                                           //                                           uart_0_s1.address
		.uart_0_s1_write                                             (mm_interconnect_0_uart_0_s1_write),                                             //                                                    .write
		.uart_0_s1_read                                              (mm_interconnect_0_uart_0_s1_read),                                              //                                                    .read
		.uart_0_s1_readdata                                          (mm_interconnect_0_uart_0_s1_readdata),                                          //                                                    .readdata
		.uart_0_s1_writedata                                         (mm_interconnect_0_uart_0_s1_writedata),                                         //                                                    .writedata
		.uart_0_s1_begintransfer                                     (mm_interconnect_0_uart_0_s1_begintransfer),                                     //                                                    .begintransfer
		.uart_0_s1_chipselect                                        (mm_interconnect_0_uart_0_s1_chipselect)                                         //                                                    .chipselect
	);

	main_system_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (nios2_fft_irq_irq)                   //    sender.irq
	);

	main_system_irq_mapper irq_mapper_001 (
		.clk           (pll_outclk0_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_001_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_sound_acquisition_irq_irq)     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                                    // reset_in0.reset
		.reset_in1      (nios2_sound_acquisition_debug_reset_request_reset), // reset_in1.reset
		.reset_in2      (nios2_fft_debug_reset_request_reset),               // reset_in2.reset
		.clk            (pll_outclk1_clk),                                   //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),                    // reset_out.reset
		.reset_req      (),                                                  // (terminated)
		.reset_req_in0  (1'b0),                                              // (terminated)
		.reset_req_in1  (1'b0),                                              // (terminated)
		.reset_req_in2  (1'b0),                                              // (terminated)
		.reset_in3      (1'b0),                                              // (terminated)
		.reset_req_in3  (1'b0),                                              // (terminated)
		.reset_in4      (1'b0),                                              // (terminated)
		.reset_req_in4  (1'b0),                                              // (terminated)
		.reset_in5      (1'b0),                                              // (terminated)
		.reset_req_in5  (1'b0),                                              // (terminated)
		.reset_in6      (1'b0),                                              // (terminated)
		.reset_req_in6  (1'b0),                                              // (terminated)
		.reset_in7      (1'b0),                                              // (terminated)
		.reset_req_in7  (1'b0),                                              // (terminated)
		.reset_in8      (1'b0),                                              // (terminated)
		.reset_req_in8  (1'b0),                                              // (terminated)
		.reset_in9      (1'b0),                                              // (terminated)
		.reset_req_in9  (1'b0),                                              // (terminated)
		.reset_in10     (1'b0),                                              // (terminated)
		.reset_req_in10 (1'b0),                                              // (terminated)
		.reset_in11     (1'b0),                                              // (terminated)
		.reset_req_in11 (1'b0),                                              // (terminated)
		.reset_in12     (1'b0),                                              // (terminated)
		.reset_req_in12 (1'b0),                                              // (terminated)
		.reset_in13     (1'b0),                                              // (terminated)
		.reset_req_in13 (1'b0),                                              // (terminated)
		.reset_in14     (1'b0),                                              // (terminated)
		.reset_req_in14 (1'b0),                                              // (terminated)
		.reset_in15     (1'b0),                                              // (terminated)
		.reset_req_in15 (1'b0)                                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                                    // reset_in0.reset
		.reset_in1      (nios2_sound_acquisition_debug_reset_request_reset), // reset_in1.reset
		.reset_in2      (nios2_fft_debug_reset_request_reset),               // reset_in2.reset
		.clk            (pll_outclk0_clk),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),                // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req),            //          .reset_req
		.reset_req_in0  (1'b0),                                              // (terminated)
		.reset_req_in1  (1'b0),                                              // (terminated)
		.reset_req_in2  (1'b0),                                              // (terminated)
		.reset_in3      (1'b0),                                              // (terminated)
		.reset_req_in3  (1'b0),                                              // (terminated)
		.reset_in4      (1'b0),                                              // (terminated)
		.reset_req_in4  (1'b0),                                              // (terminated)
		.reset_in5      (1'b0),                                              // (terminated)
		.reset_req_in5  (1'b0),                                              // (terminated)
		.reset_in6      (1'b0),                                              // (terminated)
		.reset_req_in6  (1'b0),                                              // (terminated)
		.reset_in7      (1'b0),                                              // (terminated)
		.reset_req_in7  (1'b0),                                              // (terminated)
		.reset_in8      (1'b0),                                              // (terminated)
		.reset_req_in8  (1'b0),                                              // (terminated)
		.reset_in9      (1'b0),                                              // (terminated)
		.reset_req_in9  (1'b0),                                              // (terminated)
		.reset_in10     (1'b0),                                              // (terminated)
		.reset_req_in10 (1'b0),                                              // (terminated)
		.reset_in11     (1'b0),                                              // (terminated)
		.reset_req_in11 (1'b0),                                              // (terminated)
		.reset_in12     (1'b0),                                              // (terminated)
		.reset_req_in12 (1'b0),                                              // (terminated)
		.reset_in13     (1'b0),                                              // (terminated)
		.reset_req_in13 (1'b0),                                              // (terminated)
		.reset_in14     (1'b0),                                              // (terminated)
		.reset_req_in14 (1'b0),                                              // (terminated)
		.reset_in15     (1'b0),                                              // (terminated)
		.reset_req_in15 (1'b0)                                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_fft_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_outclk0_clk),                     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                                    // reset_in0.reset
		.reset_in1      (nios2_sound_acquisition_debug_reset_request_reset), // reset_in1.reset
		.reset_in2      (nios2_fft_debug_reset_request_reset),               // reset_in2.reset
		.clk            (),                                                  //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),                // reset_out.reset
		.reset_req      (),                                                  // (terminated)
		.reset_req_in0  (1'b0),                                              // (terminated)
		.reset_req_in1  (1'b0),                                              // (terminated)
		.reset_req_in2  (1'b0),                                              // (terminated)
		.reset_in3      (1'b0),                                              // (terminated)
		.reset_req_in3  (1'b0),                                              // (terminated)
		.reset_in4      (1'b0),                                              // (terminated)
		.reset_req_in4  (1'b0),                                              // (terminated)
		.reset_in5      (1'b0),                                              // (terminated)
		.reset_req_in5  (1'b0),                                              // (terminated)
		.reset_in6      (1'b0),                                              // (terminated)
		.reset_req_in6  (1'b0),                                              // (terminated)
		.reset_in7      (1'b0),                                              // (terminated)
		.reset_req_in7  (1'b0),                                              // (terminated)
		.reset_in8      (1'b0),                                              // (terminated)
		.reset_req_in8  (1'b0),                                              // (terminated)
		.reset_in9      (1'b0),                                              // (terminated)
		.reset_req_in9  (1'b0),                                              // (terminated)
		.reset_in10     (1'b0),                                              // (terminated)
		.reset_req_in10 (1'b0),                                              // (terminated)
		.reset_in11     (1'b0),                                              // (terminated)
		.reset_req_in11 (1'b0),                                              // (terminated)
		.reset_in12     (1'b0),                                              // (terminated)
		.reset_req_in12 (1'b0),                                              // (terminated)
		.reset_in13     (1'b0),                                              // (terminated)
		.reset_req_in13 (1'b0),                                              // (terminated)
		.reset_in14     (1'b0),                                              // (terminated)
		.reset_req_in14 (1'b0),                                              // (terminated)
		.reset_in15     (1'b0),                                              // (terminated)
		.reset_req_in15 (1'b0)                                               // (terminated)
	);

endmodule
